module lab_test(
    input wire clk,
    output wire clk_o
);

assign clk_o = clk;

endmodule